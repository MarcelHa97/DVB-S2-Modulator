----------------------------------------------------------------------------------
-- Company: SeeSat e.V. (DHBW-Ravensburg Campus Friedrichshafen)
-- Engineer: Mert-Can �nl�
--          
-- Create Date: 31.01.2021 16:47:46
-- Design Name: Merger-Slice 
-- Module Name: Merger_Slicer
-- Project Name: DVB-S2
-- Target Devices: Zynq-7020
-- Tool Versions: 2020.1
-- Description: The Merger Slicer stores the UP-packets in a Datafield.
--              The length of this Datafield is depending on the FEC-Rate.
--              (see talbe 5 in DVB-S2 Standard) 
--              Only entire UPs are saved in the datafield.       
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_std.all;
 
---------------------------------------------------------------------------------------------------------------------------------------------------------------------        
entity Merger_Slicer is                                                            --The worth for KBCH is depending on the FEC-Rate(see table 5 in DVB-S2 standard)
generic( Kbch_length : integer := 14232;
         UP_Packet_Length : integer := 1024);  --1769                                      -- Length of a UP packet
port(
    clk                 : in    std_logic;                                          --Clock
    enable              : in    std_logic;                                          --Indicates that the next UP is ready 
    dataUP              : in    std_logic_vector(UP_Packet_Length downto 1);                    --Here will be stored the next UP packet from the Input-Buffer
    reset               : in    std_logic;                                          --The Stream Adaption indicates that the Frame(BBHeader_Datafield) is received; Reset "frame_ready"
    BBHeader            : in    std_logic_vector(80 downto 1);                      --BBHeader which is generated by the BBSignaling Block
    
    frame_ready         : out   std_logic;                                          --Indicates to the Stream Adaption, that the Frame is ready
    BBHeader_Datafield  : out   std_logic_vector(Kbch_length downto 1);                    --Frame / 2128
    UP_reset            : out   std_logic;                                          --Indicates that one UP is stored
   
    x_out                   : out   std_logic_vector(20 downto 0);                  --Only for Simulation
    count_out               : out   std_logic_vector(20 downto 0)                   --Only for Simulation
);
end Merger_Slicer;
--------------------------------------------------------------------------------------------------------------------------------------------------------------------- 



architecture Behavioral of Merger_Slicer is
-------------------------------------------------------------------------------------------------------------------------------
--Signals 
    signal UP_reset_s             : std_logic;
-------------------------------------------------------------------------------------------------------------------------------


begin
---------------------------------------------------------------------------------------------------------------------------------------------------------------- 
    process(enable, clk, reset)
---------------------------------------------------------------------------------------------------------------------------------------------------------------- 
 --Declaration of Variable:
    variable BBHeader_Datafield_var : std_logic_vector(2 downto 1);
    variable DataUP_var             : std_logic_vector(UP_Packet_Length downto 1);
    variable Datafield_var          : std_logic_vector(Kbch_length-80 downto 1);
    variable count                  : integer            := 0;
    variable KBCH_var               : integer            := Kbch_length;                                       --Length of the Datafield
    variable x                      : integer            := 13;  --8                                        --How often does a UP(1024) fit integer into a datafield(2128):(2128-80)/1024;
    variable enable_var             : std_logic          := '0';
    variable test_ready             : std_logic;
---------------------------------------------------------------------------------------------------------------------------------------------------------------- 
    begin 
        
        DataUP_var                                       := DataUP;                                     --store the UP in a Variable
        x_out                                            <= std_logic_vector(to_unsigned(x,21));        --Only for Simulation
        
        
        if (falling_edge(clk) and enable = '1') then            
            Datafield_var := Datafield_var(Kbch_length-80-UP_Packet_Length downto 1) & DataUP_var;
            count := count + 1;
            count_out                                     <= std_logic_vector(to_unsigned(count,21));
            UP_reset_s                                    <= '1';                                        --Indicates that one UP-Packet is stored
            frame_ready                                   <= '0';
            enable_var                                    := '0';
        end if;        
 --------------------------------------------------------------------------------------------------------------------------------       
        if (count = x) then
            enable_var                                    := '1';                                        --Indicates that Datafield is already filled with UP
        end if; 
 --------------------------------------------------------------------------------------------------------------------------------                  
        if (enable_var = '1') then      
            BBHeader_Datafield(Kbch_length-80 downto 1)           <= Datafield_var;
            BBHeader_Datafield(Kbch_length downto Kbch_length-80+1)      <= BBHeader;
            count                                          := 0;
            enable_var                                     := '0';
            frame_ready                                    <= '1';                                     --Indicates that one Frame is ready
        end if;

        if (reset = '1') then                                                                           --If reset is one, then the Frame is readed by the Stream Adaption
            frame_ready                                     <= '0';  
            Datafield_var                                   := (others => '0');                         --Reset Datafield Variable                 
        end if;
           
        if (UP_reset_s = '1') then
            UP_reset_s                                      <= '0';
        end if;   
    
    end process;
----------------------------------------------------------------------------------------------------------------------------------------------------------------
UP_reset <= UP_reset_s;


end Behavioral;






